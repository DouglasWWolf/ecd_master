
//================================================================================================
//    Date         Version     Who  Changes
// -----------------------------------------------------------------------------------------------
// 29-Sep-2022     0.1.0-rc1   DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 0;
localparam VERSION_MINOR = 1;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 1;

localparam VERSION_DAY   = 29;
localparam VERSION_MONTH = 9;
localparam VERSION_YEAR  = 2022;
