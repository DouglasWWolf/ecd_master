
//================================================================================================
//    Date         Version     Who  Changes
// -----------------------------------------------------------------------------------------------
// 29-Sep-2022     0.1.0-rc1   DWW  Initial creation
//
// 28-Oct-2022     0.2.0-rc1   DWW  Running at 40 GBit/second.  DMA byte order is fixed and
//                                  restart_manager has been added
//================================================================================================
localparam VERSION_MAJOR = 0;
localparam VERSION_MINOR = 2;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 1;

localparam VERSION_DAY   = 28;
localparam VERSION_MONTH = 10;
localparam VERSION_YEAR  = 2022;
